`timescale 1ns/1ps

module SHIFT32_TB;
	reg [31:0] D, S;
	reg LnR;
	wire [31:0] Y;
	
	SHIFT32 shift32_inst_1(.Y(Y), .D(D), .S(S), .LnR(LnR));
	
	initial begin
		D = 'b0000000000000000000000001000; S = 'b0000000000000000000000000010; LnR = 'b0;
		#5 D = 'b0000000000000000000000001000; S = 'b0000000000000000000000000010; LnR = 'b1; $write("Y =: %b\n", Y);
		#5 D = 'b0000000000000000000000001000; S = 'b0000000000000000000000000100; LnR = 'b0; $write("Y =: %b\n", Y);
		#5 D = 'b0000000000000000000000001000; S = 'b0000000000000000000000000100; LnR = 'b1; $write("Y =: %b\n", Y);
		#5 D = 'b0000000000000000000000001000; S = 'b0000000000000000000000001000; LnR = 'b0; $write("Y =: %b\n", Y);
		#5 D = 'b0000000000000000000000001000; S = 'b0000000000000000000000001000; LnR = 'b1; $write("Y =: %b\n", Y);
		#5 D = 'b0000000000000000000000001000; S = 'b0000000000000000000000010000; LnR = 'b0; $write("Y =: %b\n", Y);
		#5 D = 'b0000000000000000000000001000; S = 'b0000000000000000000000010000; LnR = 'b1; $write("Y =: %b\n", Y);
		#5 D = 'b0000000000000000000000001000; S = 'b0000000000000000000000100000; LnR = 'b1; $write("Y =: %b\n", Y);
		#5 $write("Y =: %b\n", Y);
		$stop;
	end
endmodule
